- alu ✅
- aluTest ✅
- opcode ✅
- adder ✅
- shifter ✅
- mux ✅
- in und outputs ✅

✅
🚧